module notGate(input a, output out);

    not(out,a);

endmodule